module funcao_decremente (
    input wire a,       // Primeira entrada
    input wire b,       // Segunda entrada
    output wire y       // Saída
);

    // Implementação da lógica AND
assign y = a & b;

endmodule
